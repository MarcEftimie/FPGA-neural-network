
`timescale 1ns/1ps
`default_nettype none

module perceptron_top
    (
        input wire clk_i, reset_i
    );

endmodule
