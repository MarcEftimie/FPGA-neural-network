`timescale 1ns/1ps
`default_nettype none

module perceptron_top_tb;

    parameter CLK_PERIOD_NS = 10;
    logic clk_i, logic ;
    wire out1, wire ;

    perceptron_top #(
    .HELLO(HELLO),
    .HELLO2(HELLO2))
    UUT(
        .*
    );

    always #(CLK_PERIOD_NS/2) clk_i = ~clk_i;

    initial begin
        $dumpfile("perceptron_top.fst");
        $dumpvars(0, UUT);
        clk_i = 0;
        reset_i = 1;
        repeat(1) @(negedge clk_i);
        reset_i = 0;
        $finish;
    end

endmodule
