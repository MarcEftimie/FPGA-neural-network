
`timescale 1ns/1ps
`default_nettype none

module perceptron_top
    #(
        parameter HELLO = 1;
        parameter HELLO2 = 1;
    ) (
        input wire clk_i, reset_i, btn_i,
        output logic out1, led1
    );

endmodule
